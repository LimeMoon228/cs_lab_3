module Ex2_OR(x3,x2,x1,f);
input x3,x2,x1;
output f;
assign f = ~(~(~x2 | x1 ) | ~(~x3 | ~x2) | ~(~x3 | x1) | ~(x3 |x2 |~x1 ));
endmodule
library verilog;
use verilog.vl_types.all;
entity tb_Control_Dev_Volodenkov is
end tb_Control_Dev_Volodenkov;
